module moor_s1s2_rst_asyn(
    input clk, rst, x,
    output reg [1:0]state, next_s
    );
    
endmodule